/*
=================BROUGHT TO YOU BY : TARANG SMVDU======================
***********************************************************************
INSTRUCTION => Sample Code Snippet is provided without logic with signal/port
description
-------------------------Write your own Logic-----------------------------------------------
*/
//======================================================================================

//===============
//   1) NOT GATE
//==============

module not_gate(
    input a,
    output y
);
// write logic here
endmodule
//========================================================================================

//==================
// 2) AND GATE
//==================

module and_gate(
    input a, b,
    output y
);
// write logic here
endmodule

//=======================================================================================

//==================
// 3) OR GATE
//==================

module or_gate(
    input a, b,
    output y
);
// write logic here
endmodule

//=======================================================================================

//==================
// 4) XOR GATE
//==================

module xor_gate(
    input a, b,
    output y
);
//Write your logic here
endmodule

//=======================================================================================

//==================
// 5) HALF ADDER
//==================

module half_adder(
    input a, b,
    output sum, carry
);
// write logic here
endmodule

//======================================================================================

//==================
// 6) FULL ADDER
//==================

module full_adder(
    input a, b, cin,
    output sum, cout
);
// write logic here
endmodule

//======================================================================================

//=====================
// 7) HALF SUBTRACTOR
//=====================

module half_subtractor(
    input a, b,
    output diff, borrow
);
// write logic here
endmodule

//====================================================================================

//======================
// 8) FULL SUBTRACTOR
//======================

module full_subtractor(
    input a, b, bin,
    output diff, bout
);
// write logic here
endmodule

//===================================================================================

//==========================
// 9) DECODER 2X4
//==========================

module decoder2to4(
    input a, b,
    output d0, d1, d2, d3
);
// write logic here
endmodule

//===================================================================================

//=============================
// 10) ENCODER 4x2
//=============================

module encoder4to2(
    input d0, d1, d2, d3,
    output a, b
);
// write logic here
endmodule

//=====================================================================================

//=============================
// 11) MUX 2X1
//============================

module mux2to1(
    input a, b, sel,
    output y
);
// write logic here
endmodule
//======================================================================================



//---------------------END OF SESSION 1-------------------------------------------------


